parameter imwidth=130;
parameter imheight=130;
